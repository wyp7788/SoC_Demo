module top(


);

endmodule
